module alu;
endmodule
